../tb/testbench.sv